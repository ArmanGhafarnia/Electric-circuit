** Profile: "SCHEMATIC1-p3"  [ D:\3\p3-schematic1-p3.sim ] 

** Creating circuit file "p3-schematic1-p3.sim.cir" 
** WARNING: THIS AUTOMATICALLY GENERATED FILE MAY BE OVERWRITTEN BY SUBSEQUENT SIMULATIONS

*Libraries: 
* Local Libraries :
* From [PSPICE NETLIST] section of C:\Program Files\Orcad\PSpice\PSpice.ini file:
.lib "nom.lib" 

*Analysis directives: 
.DC LIN V_V1 4 20 1 
.PROBE V(*) I(*) W(*) D(*) NOISE(*) 
.INC ".\p3-SCHEMATIC1.net" 


.END
