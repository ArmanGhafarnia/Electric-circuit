** Profile: "SCHEMATIC1-soal4"  [ d:\4\p4-SCHEMATIC1-soal4.sim ] 

** Creating circuit file "p4-SCHEMATIC1-soal4.sim.cir" 
** WARNING: THIS AUTOMATICALLY GENERATED FILE MAY BE OVERWRITTEN BY SUBSEQUENT SIMULATIONS

*Libraries: 
* Local Libraries :
* From [PSPICE NETLIST] section of C:\Program Files\Orcad\PSpice\PSpice.ini file:
.lib "nom.lib" 

*Analysis directives: 
.DC LIN V_v1 0 10 1 
.PROBE V(*) I(*) W(*) D(*) NOISE(*) 
.INC ".\p4-SCHEMATIC1.net" 


.END
