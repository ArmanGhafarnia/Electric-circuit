** Profile: "SCHEMATIC1-3c"  [ d:\3\p3-SCHEMATIC1-3c.sim ] 

** Creating circuit file "p3-SCHEMATIC1-3c.sim.cir" 
** WARNING: THIS AUTOMATICALLY GENERATED FILE MAY BE OVERWRITTEN BY SUBSEQUENT SIMULATIONS

*Libraries: 
* Local Libraries :
* From [PSPICE NETLIST] section of C:\Program Files\Orcad\PSpice\PSpice.ini file:
.lib "nom.lib" 

*Analysis directives: 
.TRAN  0 5ns 0 
.PROBE V(*) I(*) W(*) D(*) NOISE(*) 
.INC ".\p3-SCHEMATIC1.net" 


.END
