** Profile: "SCHEMATIC1-soal1-4"  [ c:\users\mahdi\desktop\sbu\elec\project\2\1\soal1-SCHEMATIC1-soal1-4.sim ] 

** Creating circuit file "soal1-SCHEMATIC1-soal1-4.sim.cir" 
** WARNING: THIS AUTOMATICALLY GENERATED FILE MAY BE OVERWRITTEN BY SUBSEQUENT SIMULATIONS

*Libraries: 
* Local Libraries :
* From [PSPICE NETLIST] section of C:\Program Files\Orcad\PSpice\PSpice.ini file:
.lib "nom.lib" 

*Analysis directives: 
.AC DEC 1 1 200
.PROBE V(*) I(*) W(*) D(*) NOISE(*) 
.INC ".\soal1-SCHEMATIC1.net" 


.END
