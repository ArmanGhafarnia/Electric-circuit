** Profile: "SCHEMATIC1-soal2-1"  [ c:\users\mahdi\desktop\sbu\elec\project\2\2\soal2-schematic1-soal2-1.sim ] 

** Creating circuit file "soal2-schematic1-soal2-1.sim.cir" 
** WARNING: THIS AUTOMATICALLY GENERATED FILE MAY BE OVERWRITTEN BY SUBSEQUENT SIMULATIONS

*Libraries: 
* Local Libraries :
* From [PSPICE NETLIST] section of C:\Program Files\Orcad\PSpice\PSpice.ini file:
.lib "nom.lib" 

*Analysis directives: 
.TRAN  0 0.5 0 
.PROBE V(*) I(*) W(*) D(*) NOISE(*) 
.INC ".\soal2-SCHEMATIC1.net" 


.END
