** Profile: "SCHEMATIC1-soal1-2"  [ D:\1-22\1-2-SCHEMATIC1-soal1-2.sim ] 

** Creating circuit file "1-2-SCHEMATIC1-soal1-2.sim.cir" 
** WARNING: THIS AUTOMATICALLY GENERATED FILE MAY BE OVERWRITTEN BY SUBSEQUENT SIMULATIONS

*Libraries: 
* Local Libraries :
* From [PSPICE NETLIST] section of C:\Program Files\Orcad\PSpice\PSpice.ini file:
.lib "nom.lib" 

*Analysis directives: 
.TRAN  0 10 0 
.PROBE V(*) I(*) W(*) D(*) NOISE(*) 
.INC ".\1-2-SCHEMATIC1.net" 


.END
